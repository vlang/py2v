@[translated]
module main

pub struct OpType {
pub mut:
	add Callable
	mul Callable
}
