@[translated]
module main

fn show() {
	// try {
	(3 / 0)
	// } catch {
	// except ZeroDivisionError:
	// NOTE: V uses Result types (!) and or{} blocks instead of exceptions
	// println('ZeroDivisionError')
	// }
}

fn main() {
	show()
}
