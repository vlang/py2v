@[translated]
module main

__global (
	num1 = 15
	num2 = 12
	sum = (num1 + num2)
)

fn main() {
	num1 = 0
	num2 = 0
	println(('Sum of {0} and {1} is {2}' /* .format(num1, num2, sum) not supported */).str())
}
