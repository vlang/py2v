@[translated]
module main

fn main_func() {
	sys.stdout.write('foobar\n')
}

fn main() {
	main_func()
}
