@[translated]
module main

fn main() {
	a := 10
	println((['hello ', ((a + 1)).str(), ' world'].join('')).str())
}
