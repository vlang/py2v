@[translated]
module main

fn main_func() {
	println('Hello, World!')
}

fn main() {
	main_func()
}
