@[translated]
module main

import math

fn main_func() {
	a := math.powi(2, 4)
	println(a.str())
}

fn main() {
	main_func()
}
