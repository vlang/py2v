@[translated]
module main

fn show() {
	// try {
	(3 / 0)
	// } catch {
	// except ZeroDivisionError:
	// NOTE: V does not have exception handling - this code is unreachable
	// println('ZeroDivisionError')
	// }
}

fn main() {
	show()
}
